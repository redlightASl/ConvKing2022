module hist_top_tb();




endmodule