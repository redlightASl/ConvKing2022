`timescale 1ns/1ps

module mobilenet_top(

);

yolo_mobilenet yolo_body(

);

endmodule
