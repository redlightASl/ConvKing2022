`timescale 1ns/1ps

module yolo_pre(

);


//get origin image



//resize



//convert to rgb888

endmodule
