`timescale 1ns/1ps

module frame_fifo_read #(
           parameter MEM_DATA_BITS = 32,
           parameter ADDR_BITS = 23,
           parameter BUSRT_BITS = 10,
           parameter FIFO_DEPTH = 256,
           parameter BURST_SIZE = 128
       )
       (
           input rst,
           input mem_clk,                     // external memory controller user interface clock
           output reg rd_burst_req,                // to external memory controller,send out a burst read request
           output reg[BUSRT_BITS - 1: 0] rd_burst_len,                // to external memory controller,data length of the burst read request, not bytes
           output reg[ADDR_BITS - 1: 0] rd_burst_addr,               // to external memory controller,base address of the burst read request
           input rd_burst_data_valid,         // from external memory controller,read request data valid
           input rd_burst_finish,             // from external memory controller,burst read finish
           input read_req,                    // data read module read request,keep '1' until read_req_ack = '1'
           output reg read_req_ack,                // data read module read request response
           output read_finish,                 // data read module read request finish
           input[ADDR_BITS - 1: 0] read_addr_0,                 // data read module read request base address 0, used when read_addr_index = 0
           input[ADDR_BITS - 1: 0] read_addr_1,                 // data read module read request base address 1, used when read_addr_index = 1
           input[ADDR_BITS - 1: 0] read_addr_2,                 // data read module read request base address 1, used when read_addr_index = 2
           input[ADDR_BITS - 1: 0] read_addr_3,                 // data read module read request base address 1, used when read_addr_index = 3
           input[1: 0] read_addr_index,             // select valid base address from read_addr_0 read_addr_1 read_addr_2 read_addr_3
           input[ADDR_BITS - 1: 0] read_len,                    // data read module read request data length
           output reg fifo_aclr,                   // to fifo asynchronous clear
           input[15: 0] wrusedw                     // from fifo write used words
       );
localparam ONE = 256'd1;                   //256 bit '1'   you can use ONE[n-1:0] for n bit '1'
localparam ZERO = 256'd0;                   //256 bit '0'
//read state machine code
localparam S_IDLE = 0;                        //idle state,waiting for frame read
localparam S_ACK = 1;                        //read request response
localparam S_WAIT = 2;
localparam S_CHECK_FIFO = 3;                        //check the FIFO status, ensure that there is enough space to burst read
localparam S_READ_BURST = 4;                        //begin a burst read
localparam S_READ_BURST_END = 5;                        //a burst read complete
localparam S_END = 6;                        //a frame of data is read to complete

reg read_req_d0;                //asynchronous read request, synchronize to 'mem_clk' clock domain,first beat
reg read_req_d1;                //second
reg read_req_d2;                //third,Why do you need 3 ? Here's the design habit
reg[ADDR_BITS - 1: 0] read_len_d0;                //asynchronous read_len(read data length), synchronize to 'mem_clk' clock domain first
reg[ADDR_BITS - 1: 0] read_len_d1;                //second
reg[ADDR_BITS - 1: 0] read_len_latch;             //lock read data length
reg[ADDR_BITS - 1: 0] read_cnt;                   //read data counter
reg[3: 0] state;                      //state machine
reg[1: 0] read_addr_index_d0;         //synchronize to 'mem_clk' clock domain first
reg[1: 0] read_addr_index_d1;         //synchronize to 'mem_clk' clock domain second
reg[15: 0] wait_cnt;
assign read_finish = (state == S_END) ? 1'b1 : 1'b0;             //read finish at state 'S_END'
always@(posedge mem_clk or posedge rst) begin
    if (rst == 1'b1) begin
        read_req_d0 <= 1'b0;
        read_req_d1 <= 1'b0;
        read_req_d2 <= 1'b0;
        read_len_d0 <= ZERO[ADDR_BITS - 1: 0];               //equivalent to read_len_d0 <= 0;
        read_len_d1 <= ZERO[ADDR_BITS - 1: 0];               //equivalent to read_len_d1 <= 0;
        read_addr_index_d0 <= 2'b00;
        read_addr_index_d1 <= 2'b00;
    end
    else begin
        read_req_d0 <= read_req;
        read_req_d1 <= read_req_d0;
        read_req_d2 <= read_req_d1;
        read_len_d0 <= read_len;
        read_len_d1 <= read_len_d0;
        read_addr_index_d0 <= read_addr_index;
        read_addr_index_d1 <= read_addr_index_d0;
    end
end


always@(posedge mem_clk or posedge rst) begin
    if (rst == 1'b1) begin
        state <= S_IDLE;
        read_len_latch <= ZERO[ADDR_BITS - 1: 0];
        rd_burst_addr <= ZERO[ADDR_BITS - 1: 0];
        rd_burst_req <= 1'b0;
        read_cnt <= ZERO[ADDR_BITS - 1: 0];
        fifo_aclr <= 1'b0;
        rd_burst_len <= ZERO[BUSRT_BITS - 1: 0];
        read_req_ack <= 1'b0;
        wait_cnt <= 16'd0;
    end
    else
    case (state)
        //idle state,waiting for read, read_req_d2 == '1' goto the 'S_ACK'
        S_IDLE: begin
            if (read_req_d2 == 1'b1) begin
                state <= S_ACK;
            end
            read_req_ack <= 1'b0;
        end
        //'S_ACK' state completes the read request response, the FIFO reset, the address latch, and the data length latch
        S_ACK: begin
            if (read_req_d2 == 1'b0) begin
                state <= S_WAIT;
                wait_cnt <= 16'd0;
                fifo_aclr <= 1'b0;
                read_req_ack <= 1'b0;
            end
            else begin
                //read request response
                read_req_ack <= 1'b1;
                //FIFO reset
                fifo_aclr <= 1'b1;
                //select valid base address from read_addr_0 read_addr_1 read_addr_2 read_addr_3
                if (read_addr_index_d1 == 2'd0)
                    rd_burst_addr <= read_addr_0;
                else if (read_addr_index_d1 == 2'd1)
                    rd_burst_addr <= read_addr_1;
                else if (read_addr_index_d1 == 2'd2)
                    rd_burst_addr <= read_addr_2;
                else if (read_addr_index_d1 == 2'd3)
                    rd_burst_addr <= read_addr_3;
                //latch data length
                read_len_latch <= read_len_d1;
            end
            //read data counter reset, read_cnt <= 0;
            read_cnt <= ZERO[ADDR_BITS - 1: 0];
        end
        S_WAIT: begin
            if (wait_cnt >= 16'd200) begin
                state <= S_CHECK_FIFO;
            end
            else begin
                wait_cnt <= wait_cnt + 16'd1;
            end
        end
        S_CHECK_FIFO: begin
            //if there is a read request at this time, enter the 'S_ACK' state
            if (read_req_d2 == 1'b1) begin
                state <= S_ACK;
            end
            //if the FIFO space is a burst read request, goto burst read state
            else if (wrusedw < (FIFO_DEPTH - BURST_SIZE - 2)) begin
                state <= S_READ_BURST;
                rd_burst_len <= BURST_SIZE[BUSRT_BITS - 1: 0];
                rd_burst_req <= 1'b1;
            end
        end

        S_READ_BURST: begin
            if (rd_burst_data_valid)
                rd_burst_req <= 1'b0;
            //burst finish
            if (rd_burst_finish == 1'b1) begin
                state <= S_READ_BURST_END;
                //read counter + burst length
                read_cnt <= read_cnt + BURST_SIZE[ADDR_BITS - 1: 0];
                //the next burst read address is generated
                rd_burst_addr <= rd_burst_addr + BURST_SIZE[ADDR_BITS - 1: 0];
            end
        end
        S_READ_BURST_END: begin
            //if there is a read request at this time, enter the 'S_ACK' state
            if (read_req_d2 == 1'b1) begin
                state <= S_ACK;
            end
            //if the read counter value is less than the frame length, continue read,
            //otherwise the read is complete
            else if (read_cnt < read_len_latch) begin
                state <= S_CHECK_FIFO;
            end
            else begin
                state <= S_END;
            end
        end
        S_END: begin
            state <= S_IDLE;
        end
        default:
            state <= S_IDLE;
    endcase
end
endmodule
