`timescale 1ns/1ps

module mobilenet_invers(

       );


yolo_cbl cbl_layer_1
(
);

endmodule
