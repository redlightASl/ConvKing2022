`timescale 1ns/1ps

module yolo_mobilenet(
    
);


mobilenet_invers mobilenet_invers_layer_1(

);

endmodule